`ifndef SPI_PKG
`define SPI_PKG

package spi_pkg;
	`include "transaction.sv"
	`include "generator.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "scoreboard.sv"
	`include "environment.sv"
endpackage

`endif